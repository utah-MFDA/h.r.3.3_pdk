

** Capacitor test case

*.ic v(out)=0
**.verilog "capacitor.va"

V1 1 0 PWL(0s 0V 5ms 0V 5.001ms 5V 10ms 5V)
R1 1 2 5k
*

Vp 2 3 0V
Ymembrane_cap_20pxV 3 0 1u

.tran 0.01ms 10ms

*.print tran V(2) V(1)
.print tran I(Vp)

.end