

*Vpp 1  0 PWL(0s 0V 3s 20V)
Vpp  6  0 5V

Vcc  11 0 5V

Vpn1 101 0 0V
*PWL(0s 0V 2s 0V 3s 16V 5s 16V)

Vpn2 102 0 0V
*PWL(0s 16V 3s 16V 4s 0V 5s 0V)

Yserpentine_100px_0  serp1 0 21 11 12

* probe
Vpr2 21 22 0V

Yserpentine_100px_0   serpE 22 31 11 13

* probe
Vpr1 31 32 0V

Yserpentine_100px_0  serp2 4 32 11 14

Yserpentine_100px_0  serp3 6 5 11 16
Yvalve_20px_1        valv1 5 4 11 15 101 0

Yvalve_20px_1        valv2 4 7 11 17 102 0
Yserpentine_100px_0  serp4 7 0 11 18


.tran 100ms 5s
.print tran V(22) V(31) I(Vpr1) I(Vpr2)
.end