MACRO diffmix_25px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN diffmix_25px_0 0 0 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN a_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END a_fluid
  PIN b_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END b_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 53 53 67 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 60 60 ;
    LAYER met2 ;
      RECT 30 30 60 60 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END diffmix_25px_0
