*Test of the pump object

YPressurePump prpump 1 0 pressure=100k

YChannel chan1 1 0 0 0 length=100m

.tran 1m 10m
.print tran V(1)
.end
