VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO serpentine_100px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_100px_0 0 0 ;
  SIZE 180 BY 180 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 143 23 157 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 37 37 143 143 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_100px_0
 
MACRO serpentine_150px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_150px_0 0 0 ;
  SIZE 240 BY 240 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203 23 217 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 210 210 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_150px_0
 
MACRO serpentine_200_100px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_200_100px_0 0 0 ;
  SIZE 300 BY 180 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 263 23 277 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 270 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_200_100px_0

MACRO serpentine_200px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_200px_0 0 0 ;
  SIZE 300 BY 300 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 263 23 277 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 270 270 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_200px_0
 
MACRO serpentine_200px_3
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_200px_0 0 0 ;
  SIZE 300 BY 300 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 23 23 37 37 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 30 0 270 300 ;
    LAYER met3 ;
      RECT 60 0 270 300 ;
    LAYER met4 ;
      RECT 60 0 270 300 ;
    LAYER met5 ;
      RECT 30 0 270 300 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_200px_3

MACRO serpentine_300px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 420 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 383 23 397 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 360 390 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_0

MACRO serpentine_300px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 420 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53 23 67 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23 23 37 37 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 60 0 390 420 ;
    LAYER met3 ;
      RECT 60 0 390 420 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_1
 
MACRO serpentine_300px_2
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 450 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 413 23 427 37 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 30 0 390 420 ;
    LAYER met3 ;
      RECT 60 0 390 420 ;
    LAYER met4 ;
      RECT 60 0 420 420 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_2
 
MACRO serpentine_300px_3
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 420 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53 23 67 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 23 23 37 37 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 60 0 420 420 ;
    LAYER met3 ;
      RECT 60 0 420 420 ;
    LAYER met4 ;
      RECT 60 0 420 420 ;
    LAYER met5 ;
      RECT 30 0 420 420 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_3
 
MACRO serpentine_300px_4
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 450 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met6 ;
        RECT 413 23 427 37 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 30 0 390 420 ;
    LAYER met3 ;
      RECT 60 0 390 420 ;
    LAYER met4 ;
      RECT 60 0 420 420 ;
    LAYER met5 ;
      RECT 60 0 420 420 ;
    LAYER met6 ;
      RECT 60 0 420 420 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_4
 
MACRO serpentine_50px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_50px_0 0 0 ;
  SIZE 120 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 83 23 97 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 90 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_50px_0
 
MACRO serpentine_75px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_75px_0 0 0 ;
  SIZE 150 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 113 23 127 37 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 120 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_75px_0
MACRO diffmix_25px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN diffmix_25px_0 0 0 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN a_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END a_fluid
  PIN b_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 23 37 37 ;
    END
  END b_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 53 53 67 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 37 37 53 53 ;
    LAYER met2 ;
      RECT 37 37 53 53 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END diffmix_25px_0
 
MACRO mixer_sw_test
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN mixer_sw_test 0 0 ;
  SIZE 210 BY 260 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN a_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END a_fluid
  PIN b_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.5 29.5 164.5 30.5 ;
    END
  END b_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.5 229.5 100.5 230.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 230 ;
    LAYER met2 ;
      RECT 30 30 180 230 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END mixer_sw_test

MACRO directional_res_1000nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN directional_res_1000nl 0 0 ;
  SIZE 245 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met8 ;
        RECT 23 66 37 80 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 208 66 222 80 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 20 215 130 ;
    LAYER met2 ;
      RECT 30 20 215 130 ;
    LAYER met3 ;
      RECT 30 20 215 130 ;
    LAYER met4 ;
      RECT 30 20 215 130 ;
    LAYER met5 ;
      RECT 30 20 215 130 ;
    LAYER met6 ;
      RECT 30 20 215 130 ;
    LAYER met7 ;
      RECT 30 20 215 130 ;
    LAYER met8 ;
      RECT 30 20 215 130 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END directional_res_1000nl

MACRO directional_res_400nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN directional_res_400nl 0 0 ;
  SIZE 210 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 120 ;
    LAYER met2 ;
      RECT 30 30 180 120 ;
    LAYER met3 ;
      RECT 30 30 180 120 ;
    LAYER met4 ;
      RECT 30 30 180 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END directional_res_400nl

MACRO directional_res_600nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN directional_res_600nl 0 0 ;
  SIZE 210 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met6 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 120 ;
    LAYER met2 ;
      RECT 30 30 180 120 ;
    LAYER met3 ;
      RECT 30 30 180 120 ;
    LAYER met4 ;
      RECT 30 30 180 120 ;
    LAYER met5 ;
      RECT 30 30 180 120 ;
    LAYER met6 ;
      RECT 30 30 180 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END directional_res_600nl

MACRO directional_res_800nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN directional_res_800nl 0 0 ;
  SIZE 210 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met8 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 120 ;
    LAYER met2 ;
      RECT 30 30 180 120 ;
    LAYER met3 ;
      RECT 30 30 180 120 ;
    LAYER met4 ;
      RECT 30 30 180 120 ;
    LAYER met5 ;
      RECT 30 30 180 120 ;
    LAYER met6 ;
      RECT 30 30 180 120 ;
    LAYER met7 ;
      RECT 30 30 180 120 ;
    LAYER met8 ;
      RECT 30 30 180 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END directional_res_800nl

MACRO inline_res_100nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN inline_res_100nl 0 0 ;
  SIZE 240 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203 53 217 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 210 90 ;
    LAYER met2 ;
      RECT 30 30 210 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END inline_res_100nl

MACRO inline_res_40nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN inline_res_40nl 0 0 ;
  SIZE 210 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 90 ;
    LAYER met2 ;
      RECT 30 30 180 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END inline_res_40nl

MACRO inline_res_60nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN inline_res_60nl 0 0 ;
  SIZE 180 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 143 53 157 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 150 90 ;
    LAYER met2 ;
      RECT 30 30 150 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END inline_res_60nl

MACRO inline_res_80nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN inline_res_80nl 0 0 ;
  SIZE 210 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 90 ;
    LAYER met2 ;
      RECT 30 30 180 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END inline_res_80nl

MACRO valve_40px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_40px_1 0 0 ;
  SIZE 180 BY 180 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 89.5 30.5 90.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 149.5 89.5 150.5 90.5 ;
    END
  END out_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 149.5 90.5 150.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 30 150 150 ;
    LAYER met2 ;
      RECT 30 30 150 150 ;
    LAYER met3 ;
      RECT 30 30 150 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_40px_1

MACRO valve_80px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_80px_1 0 0 ;
  SIZE 190 BY 190 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 89.5 30.5 90.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 149.5 89.5 150.5 90.5 ;
    END
  END out_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 149.5 90.5 150.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 30 150 150 ;
    LAYER met2 ;
      RECT 30 30 150 150 ;
    LAYER met3 ;
      RECT 30 30 150 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_80px_1

MACRO valve_80px_4way_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_80px_4way_0 0 0 ;
  SIZE 190 BY 190 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN a_fluid
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 89.5 30.5 90.5 ;
    END
  END a_fluid
  PIN b_fluid
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 149.5 89.5 150.5 90.5 ;
    END
  END b_fluid
  PIN c_fluid
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END c_fluid
  PIN d_fluid
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 89.5 149.5 90.5 150.5 ;
    END
  END d_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 59.5 90.5 60.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 119.5 90.5 120.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 30 150 150 ;
    LAYER met2 ;
      RECT 30 30 150 150 ;
    LAYER met3 ;
      RECT 60 60 120 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_80px_4way_0

MACRO pump_20_40_20px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_20_40_20px_0 0 0 ;
  SIZE 320 BY 165 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN fluid_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 89.5 30.5 90.5 ;
    END
  END fluid_in
  PIN fluid_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 299.5 89.5 300.5 90.5 ;
    END
  END fluid_out
  PIN a_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 149.5 90.5 150.5 ;
    END
  END a_out_air
  PIN b_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.5 149.5 165.5 150.5 ;
    END
  END b_out_air
  PIN c_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.5 149.5 240.5 150.5 ;
    END
  END c_out_air
  PIN a_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END a_in_air
  PIN b_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.5 29.5 165.5 30.5 ;
    END
  END b_in_air
  PIN c_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 239.5 29.5 240.5 30.5 ;
    END
  END c_in_air
  OBS
    LAYER met1 ;
      RECT 30 30 300 150 ;
    LAYER met2 ;
      RECT 30 30 300 150 ;
    LAYER met3 ;
      RECT 30 30 300 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_20_40_20px_0

MACRO pump_20px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_20px_0 0 0 ;
  SIZE 300 BY 130 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN fluid_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 64.5 30.5 65.5 ;
    END
  END fluid_in
  PIN fluid_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.5 64.5 270.5 65.5 ;
    END
  END fluid_out
  PIN air_out_a
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.5 99.5 80.5 100.5 ;
    END
  END air_out_a
  PIN air_out_b
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 99.5 150.5 100.5 ;
    END
  END air_out_b
  PIN air_out_c
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.5 99.5 220.5 100.5 ;
    END
  END air_out_c
  PIN air_in_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.5 29.5 80.5 30.5 ;
    END
  END air_in_a
  PIN air_in_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 29.5 150.5 30.5 ;
    END
  END air_in_b
  PIN air_in_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.5 29.5 220.5 30.5 ;
    END
  END air_in_c
  OBS
    LAYER met1 ;
      RECT 30 30 270 100 ;
    LAYER met2 ;
      RECT 30 30 270 100 ;
    LAYER met3 ;
      RECT 30 30 270 100 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_20px_0

MACRO pump_40px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_40px_0 0 0 ;
  SIZE 290 BY 135 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 59.5 30.5 60.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.5 59.5 270.5 60.5 ;
    END
  END out_fluid
  PIN a_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END a_in_air
  PIN a_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 89.5 90.5 90.5 ;
    END
  END a_out_air
  PIN b_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 29.5 150.5 30.5 ;
    END
  END b_in_air
  PIN b_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 89.5 150.5 90.5 ;
    END
  END b_out_air
  PIN c_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.5 29.5 210.5 30.5 ;
    END
  END c_in_air
  PIN c_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.5 89.5 210.5 90.5 ;
    END
  END c_out_air
  OBS
    LAYER met1 ;
      RECT 30 30 270 90 ;
    LAYER met2 ;
      RECT 30 30 270 90 ;
    LAYER met3 ;
      RECT 30 30 270 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_40px_0

MACRO optical_measure_100_5ch
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN optical_measure_100_5ch 0 0 ;
  SIZE 360 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 323 53 337 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 330 90 ;
    LAYER met2 ;
      RECT 30 30 330 90 ;
    LAYER met3 ;
      RECT 40 30 320 90 ;
    LAYER met4 ;
      RECT 30 30 330 90 ;
    LAYER met5 ;
      RECT 40 30 320 90 ;
    LAYER met6 ;
      RECT 30 30 330 90 ;
    LAYER met7 ;
      RECT 30 30 330 90 ;
    LAYER met8 ;
      RECT 30 30 330 90 ;
    LAYER met9 ;
      RECT 30 30 330 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END optical_measure_100_5ch

MACRO optical_measure_300_5ch
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN optical_measure_300_5ch 0 0 ;
  SIZE 600 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23 68 37 82 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 563 68 577 82 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 570 120 ;
    LAYER met2 ;
      RECT 30 30 570 120 ;
    LAYER met3 ;
      RECT 40 30 560 120 ;
    LAYER met4 ;
      RECT 30 30 570 120 ;
    LAYER met5 ;
      RECT 40 30 560 120 ;
    LAYER met6 ;
      RECT 30 30 570 120 ;
    LAYER met7 ;
      RECT 30 30 570 120 ;
    LAYER met8 ;
      RECT 30 30 570 120 ;
    LAYER met9 ;
      RECT 30 30 570 120 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END optical_measure_300_5ch

MACRO pinhole_325px_0
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_0 ;
  SIZE 330 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 310 60 330 80 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 60 20 80 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 20 0 310 140 ;
    LAYER met2 ;
      RECT 20 0 310 140 ;
    LAYER met3 ;
      RECT 20 0 310 140 ;
    LAYER met4 ;
      RECT 20 0 310 140 ;
    LAYER met5 ;
      RECT 20 0 310 140 ;
    LAYER met6 ;
      RECT 20 0 310 140 ;
    LAYER met7 ;
      RECT 20 0 310 140 ;
    LAYER met8 ;
      RECT 20 0 310 140 ;
    LAYER met9 ;
      RECT 20 0 310 140 ;
  END
END pinhole_325px_0
END LIBRARY
