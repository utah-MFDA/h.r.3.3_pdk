* serpentine 100 test


YPressurePump pr1  1  2   pressure=100k chemConcentration=100m

Ychannel serp1 11 1 3 2 length=10m
Ychannel serp2 0 11 4 3 length=10m
*YOutput  out   4
*VCC 4 0 0V

*.preprocess addresistors nodcpath 1G
*.preprocess addresistors oneterminal 1G

.tran 1m 10m
.print tran V(3) V(11) 
*I(vcc)
.end
