################################## FUNCTIONAL ##################################



################################### TESTING ####################################

MACRO valve_20px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_20px_1 0 0 ;
  SIZE 120 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 59.5 30.5 60.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 89.5 59.5 90.5 60.5 ;
    END
  END out_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.5 29.5 60.5 30.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.5 89.5 60.5 90.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 30 90 90 ;
    LAYER met2 ;
      RECT 30 30 90 90 ;
    LAYER met3 ;
      RECT 30 30 90 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_20px_1