VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

################################## FUNCTIONAL ##################################

MACRO serpentine_50px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_50px_0 0 0 ;
  SIZE 120 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 90 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_50px_0

MACRO serpentine_100px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_100px_0 0 0 ;
  SIZE 180 BY 180 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 149.5 29.5 150.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 150 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_100px_0

MACRO serpentine_150px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_150px_0 0 0 ;
  SIZE 240 BY 240 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 209.5 29.5 210.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 210 210 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_150px_0

MACRO serpentine_200px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_200px_0 0 0 ;
  SIZE 300 BY 300 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.5 29.5 270.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 270 270 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_200px_0

MACRO serpentine_300px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 420 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 389.5 29.5 390.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 360 390 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_0








