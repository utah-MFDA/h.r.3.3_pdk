
vsi 1  0 0V

vsp 31 0 PWL(0s 0V 1ms 0kV 2ms 69kV 100ms 69kV)

r1 1 2 3e12
r2 4 0 3e12

*module valve_fl_20px_1_V2(fl_in, fl_out,  pn_in);
Yvalve_fl_20px_1_V1 valv1 2 3 31 threshold_pressure_kPa=66e3

vp1 3 4 0V

.tran 0.01ms 20ms 0s 1ms
.print tran I(vp1) V(31)
.end
