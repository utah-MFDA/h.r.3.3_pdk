

vs_f 1  0 5V
vs_p1 11 0 PWL(0s 105kV 3 105kV 3.1 0kV   12 0kV   12.1   105kV 20 105kV)
vs_p2 12 0 PWL(0s 0V    6 0v    6.1 105kV 15 105kV 15.1   0V    20 0kV)
vs_p3 13 0 PWL(0s 105kV 9 105kV 9.1 0kV   18 0kV   18.1   105kV 20 105kV)

r1 1 2 1k
r2 5 0 1k


Yvalve_20px_1_V        valv1 3 31 11 0  
Ymembrane_cap_20pxV_Pn mem1  31 12
Yvalve_20px_1_V        valv2 31 4 13 0  

vp1 3 2 0V
vp2 5 4 0V 

.tran 0.01 20s
.print tran I(vp1) I(vp2) V(11) V(12) V(13)
.end
