MACRO interconnect_8x4
  CLASS PAD ;
  SIZE 650 BY 290 ;
  ORIGIN 0 0 ;
  PIN connection_0_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 0 20 20 ;
    END
  END connection_0_0
  PIN pad_0_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 0 20 20 ;
    END
  END pad_0_0
  PIN connection_0_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 90 20 110 ;
    END
  END connection_0_1
  PIN pad_0_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 90 20 110 ;
    END
  END pad_0_1
  PIN connection_0_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 180 20 200 ;
    END
  END connection_0_2
  PIN pad_0_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 180 20 200 ;
    END
  END pad_0_2
  PIN connection_0_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 270 20 290 ;
    END
  END connection_0_3
  PIN pad_0_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 270 20 290 ;
    END
  END pad_0_3
  PIN connection_1_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 0 110 20 ;
    END
  END connection_1_0
  PIN pad_1_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 0 110 20 ;
    END
  END pad_1_0
  PIN connection_1_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 90 110 110 ;
    END
  END connection_1_1
  PIN pad_1_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 90 110 110 ;
    END
  END pad_1_1
  PIN connection_1_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 180 110 200 ;
    END
  END connection_1_2
  PIN pad_1_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 180 110 200 ;
    END
  END pad_1_2
  PIN connection_1_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 270 110 290 ;
    END
  END connection_1_3
  PIN pad_1_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 270 110 290 ;
    END
  END pad_1_3
  PIN connection_2_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 0 200 20 ;
    END
  END connection_2_0
  PIN pad_2_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 0 200 20 ;
    END
  END pad_2_0
  PIN connection_2_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 90 200 110 ;
    END
  END connection_2_1
  PIN pad_2_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 90 200 110 ;
    END
  END pad_2_1
  PIN connection_2_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 180 200 200 ;
    END
  END connection_2_2
  PIN pad_2_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 180 200 200 ;
    END
  END pad_2_2
  PIN connection_2_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 270 200 290 ;
    END
  END connection_2_3
  PIN pad_2_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 270 200 290 ;
    END
  END pad_2_3
  PIN connection_3_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 0 290 20 ;
    END
  END connection_3_0
  PIN pad_3_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 0 290 20 ;
    END
  END pad_3_0
  PIN connection_3_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 90 290 110 ;
    END
  END connection_3_1
  PIN pad_3_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 90 290 110 ;
    END
  END pad_3_1
  PIN connection_3_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 180 290 200 ;
    END
  END connection_3_2
  PIN pad_3_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 180 290 200 ;
    END
  END pad_3_2
  PIN connection_3_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 270 290 290 ;
    END
  END connection_3_3
  PIN pad_3_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 270 290 290 ;
    END
  END pad_3_3
  PIN connection_4_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 0 380 20 ;
    END
  END connection_4_0
  PIN pad_4_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 0 380 20 ;
    END
  END pad_4_0
  PIN connection_4_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 90 380 110 ;
    END
  END connection_4_1
  PIN pad_4_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 90 380 110 ;
    END
  END pad_4_1
  PIN connection_4_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 180 380 200 ;
    END
  END connection_4_2
  PIN pad_4_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 180 380 200 ;
    END
  END pad_4_2
  PIN connection_4_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 270 380 290 ;
    END
  END connection_4_3
  PIN pad_4_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 270 380 290 ;
    END
  END pad_4_3
  PIN connection_5_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 0 470 20 ;
    END
  END connection_5_0
  PIN pad_5_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 0 470 20 ;
    END
  END pad_5_0
  PIN connection_5_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 90 470 110 ;
    END
  END connection_5_1
  PIN pad_5_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 90 470 110 ;
    END
  END pad_5_1
  PIN connection_5_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 180 470 200 ;
    END
  END connection_5_2
  PIN pad_5_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 180 470 200 ;
    END
  END pad_5_2
  PIN connection_5_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 270 470 290 ;
    END
  END connection_5_3
  PIN pad_5_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 270 470 290 ;
    END
  END pad_5_3
  PIN connection_6_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 0 560 20 ;
    END
  END connection_6_0
  PIN pad_6_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 0 560 20 ;
    END
  END pad_6_0
  PIN connection_6_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 90 560 110 ;
    END
  END connection_6_1
  PIN pad_6_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 90 560 110 ;
    END
  END pad_6_1
  PIN connection_6_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 180 560 200 ;
    END
  END connection_6_2
  PIN pad_6_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 180 560 200 ;
    END
  END pad_6_2
  PIN connection_6_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 270 560 290 ;
    END
  END connection_6_3
  PIN pad_6_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 270 560 290 ;
    END
  END pad_6_3
  PIN connection_7_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 0 650 20 ;
    END
  END connection_7_0
  PIN pad_7_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 0 650 20 ;
    END
  END pad_7_0
  PIN connection_7_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 90 650 110 ;
    END
  END connection_7_1
  PIN pad_7_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 90 650 110 ;
    END
  END pad_7_1
  PIN connection_7_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 180 650 200 ;
    END
  END connection_7_2
  PIN pad_7_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 180 650 200 ;
    END
  END pad_7_2
  PIN connection_7_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 270 650 290 ;
    END
  END connection_7_3
  PIN pad_7_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 270 650 290 ;
    END
  END pad_7_3
END interconnect_8x4
