
MACRO inline_res_80nl
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN inline_res_80nl 0 0 ;
  SIZE 210 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173 53 187 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 180 90 ;
    LAYER met2 ;
      RECT 30 30 180 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END inline_res_80nl
