
MACRO pump_20px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_20px_0 0 0 ;
  SIZE 300 BY 150 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN fluid_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 62.5 30.5 63.5 ;
    END
  END fluid_in
  PIN fluid_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269 62.5 270.5 63.5 ;
    END
  END fluid_out
  PIN air_out_a
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.5 99.5 78.5 100.5 ;
    END
  END air_out_a
  PIN air_out_b
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.5 99.5 148.5 100.5 ;
    END
  END air_out_b
  PIN air_out_c
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.5 99.5 218.5 100.5 ;
    END
  END air_out_c
  PIN air_in_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.5 29.5 78.5 30.5 ;
    END
  END air_in_a
  PIN air_in_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.5 29.5 148.5 30.5 ;
    END
  END air_in_b
  PIN air_in_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.5 29.5 218.5 30.5 ;
    END
  END air_in_c
  OBS
    LAYER met1 ;
      RECT 30 30 280 110 ;
    LAYER met2 ;
      RECT 30 30 280 110 ;
    LAYER met3 ;
      RECT 30 30 280 110 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_20px_0
