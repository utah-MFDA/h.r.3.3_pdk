* one stop valve per device

vs_f 1  0 0V

vs_p1 11 0 PULSE(69kV 0kV   0.56   5m 5m 60m  300m)
vs_p2 12 0 PULSE(69kV 0kV   0.561  5m 5m 180m 300m)
vs_p3 13 0 PULSE(69kV 0kV   0.68   5m 5m 120m 300m)

r1 1 2 1e12
r2 5 0 1e12


Yvalve_sw_20px_1_V              valv1 3  31 11 0 threshold_pressure_kPa=60e3 
Ymembrane_cap_20pxV_nlin_5_1 mem1  31 12 mem_r=504e-6 fl_ch_h=60e-6
Yvalve_sw_20px_1_V              valv2 31 4 13 0 threshold_pressure_kPa=60e3 

vp1 2 3 0V
vp2 4 5 0V 

.tran 0.01ms 2.1s 0.4s 0.1ms
.print tran I(vp1) I(vp2) V(11) V(12) V(13)
.end
