
vsi 1  0 0V

vsp 31 0 PWL(0s 0V 1ms 0kV 2ms 69kV 100ms 69kV)

r1 1 2 1e11
r2 4 0 1e11

*module valve_fl_20px_1_V2(fl_in, fl_out,  pn_in);

Yvalve_sw_20px_1_V           valv1 2 3 31 0 threshold_pressure_kPa=68e3
Ymembrane_cap_20pxV_nlin_3_1 mem1  3 31 mem_r=540e-6 fl_ch_h=60e-6

vp1 3 4 0V

.tran 0.01ms 20ms 0s 1ms
.print tran I(vp1) I(vsi) V(31)
.end
