

vs1  1  0 10k
vsc1 11 0 0

Ychannel ch1 1 2 11 12 length=10m
Ychannel ch2 2 0 12 13 length=10m

.tran 0.1ms 1
.print tran V(1) V(11) I(vs1)
.end

