// q_in, flow in, l, length, r, radius
module circular_channel (q_in, l, r);
