
.options linsol type=klu

vs 1 0 PWL(0s 0V 3ms 0V 3.001ms 56e3V 6.0ms 56e3V 6.001ms -56e3V 10ms -56e3V)
r1 0 11 1k
r2 13 0 1k
Ymembrane_cap_20pxV_nlin mem1 2 1 


* probe sources
vp1 11 2 0V
vp2 2 13 0V

.tran 0.001ms 10ms
*.option post=2
.print tran I(vp2) I(vp1) I(vs) V(1) V(2)
.end
