
MACRO valve_80px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_80px_1 0 0 ;
  SIZE 190 BY 190 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 89.5 30.5 90.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 149.5 89.5 150.5 90.5 ;
    END
  END out_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 29.5 90.5 30.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 149.5 90.5 150.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 30 150 150 ;
    LAYER met2 ;
      RECT 30 30 150 150 ;
    LAYER met3 ;
      RECT 30 30 150 150 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_80px_1
