

YPressurePump prPump1 1 0   pressure=100k
YPressurePump prPump2 11 0 pressure=100k

Yserpentine_100px_0 serp1 1 3 0 0
Yserpentine_100px_0 serp2 11 13 0 0

Ydiffmix_25px_0_fl mix1 3 13 5 

Yserpentine_100px_0 serp3 5 0 0 0


.tran 1m 10m 
.print tran V(1)
.end
