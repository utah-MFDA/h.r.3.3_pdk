

vs_f 1  0 5V
vs_p 11 0 PWL(0s 0V 3 0v 6 105kV 10 105kV)

r1 1 2 1k
r2 5 0 1k
*r3 11 12 1k
*r4 13 0 1M

*Yvalve_20px_1_V        valv1 3 31 11 0
r5 3 31 1.418e6
Ymembrane_cap_20pxV_Pn mem1  31 11
*Yvalve_20px_1_V        valv2 31 4 11 0  
r6 31 4 1.418e6

vp1 2 3 0V
vp2 4 5 0V 

.tran 0.01 10s
.print tran I(vp1) I(vp2)
.end