*A simple rectangular channel

.hdl ./../../RectangularChannel.va
.options post=1
X1 1 0 RectangularChannel
VS 1 0 1
.dc VS 0 10 1
.end
