

** Capacitor test case

*.ic v(out)=0
**.verilog "capacitor.va"

V1 1 0 sin( 0 2.5 20meg)
R1 1 2 5000k
R2 2 0 1000k
*
Ymembrane_cap_20pxV 2 0 1000u
*2 0 C=1000u
*
**YVLG_capacitor 0 2 capacitor
.tran 0.1n 0.5u

.print tran V(2) V(1)

.end