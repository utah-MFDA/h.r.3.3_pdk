* serpentine 100 test


YPressurePump pr1  1  2   pressure=100k chemConcentration=100m

Ychannel_flow serp1 1 11 length=10m
Ychannel_flow serp2 11 0 length=10m

*YOutput  out   4
*VCC 4 0 0V

*.preprocess addresistors nodcpath 1G
*.preprocess addresistors oneterminal 1G

.tran 1m 10m
.print tran V(11) 
*I(vcc)
.end
