

vs 1 0 5v


YOutput o1 1 0

.tran 0.1m 1m
.print tran V(1)
.end


