

vs 1 0 PWL(0s 0V 5ms 0V 5.001ms 15V 10ms 15V)
r1 1 2 1k
*c1 3 0 1uF
Ymembrane_cap_20pxV mem1 3 0
*cap=1u

vp 2 3 0V

.tran 0.01ms 10ms
*.option post=2
.print tran I(vs) I(vp) V(3) V(1)
.end