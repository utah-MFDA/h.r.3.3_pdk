
vsi 1  0 0V

vsp 31 0 PWL(0s 0V 1ms 0kV 2ms 69kV 100ms 69kV)

r1 1 2 1e12
r2 4 0 1e12

*module valve_fl_20px_1_V2(fl_in, fl_out,  pn_in);
Yvalve_fl_20px_1_V3_m5 valv1 2 3 31 mem_r=540e-6 fl_ch_h=60e-6
*threshold_pressure_kPa=60e3

vp1 3 4 0V

.tran 0.01ms 10ms 0s 1ms
.print tran I(vp1) I(vsi) V(31)
.end
