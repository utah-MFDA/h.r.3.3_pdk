VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO interconnect
  CLASS COVER BUMP ;
  SIZE 40 BY 40 ;
  ORIGIN 0 0 ;
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 0 40 40 ;
    END
  END pad
END interconnect

MACRO interconnect_8x4
  CLASS PAD ;
  SIZE 650 BY 290 ;
  ORIGIN 0 0 ;
  PIN connection_0_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 0 20 20 ;
    END
  END connection_0_0
  PIN pad_0_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 0 20 20 ;
    END
  END pad_0_0
  PIN connection_0_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 90 20 110 ;
    END
  END connection_0_1
  PIN pad_0_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 90 20 110 ;
    END
  END pad_0_1
  PIN connection_0_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 180 20 200 ;
    END
  END connection_0_2
  PIN pad_0_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 180 20 200 ;
    END
  END pad_0_2
  PIN connection_0_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 270 20 290 ;
    END
  END connection_0_3
  PIN pad_0_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 270 20 290 ;
    END
  END pad_0_3
  PIN connection_1_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 0 110 20 ;
    END
  END connection_1_0
  PIN pad_1_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 90 0 110 20 ;
    END
  END pad_1_0
  PIN connection_1_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 90 110 110 ;
    END
  END connection_1_1
  PIN pad_1_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 90 90 110 110 ;
    END
  END pad_1_1
  PIN connection_1_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 180 110 200 ;
    END
  END connection_1_2
  PIN pad_1_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 90 180 110 200 ;
    END
  END pad_1_2
  PIN connection_1_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 90 270 110 290 ;
    END
  END connection_1_3
  PIN pad_1_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 90 270 110 290 ;
    END
  END pad_1_3
  PIN connection_2_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 0 200 20 ;
    END
  END connection_2_0
  PIN pad_2_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 180 0 200 20 ;
    END
  END pad_2_0
  PIN connection_2_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 90 200 110 ;
    END
  END connection_2_1
  PIN pad_2_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 180 90 200 110 ;
    END
  END pad_2_1
  PIN connection_2_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 180 200 200 ;
    END
  END connection_2_2
  PIN pad_2_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 180 180 200 200 ;
    END
  END pad_2_2
  PIN connection_2_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 180 270 200 290 ;
    END
  END connection_2_3
  PIN pad_2_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 180 270 200 290 ;
    END
  END pad_2_3
  PIN connection_3_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 0 290 20 ;
    END
  END connection_3_0
  PIN pad_3_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 270 0 290 20 ;
    END
  END pad_3_0
  PIN connection_3_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 90 290 110 ;
    END
  END connection_3_1
  PIN pad_3_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 270 90 290 110 ;
    END
  END pad_3_1
  PIN connection_3_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 180 290 200 ;
    END
  END connection_3_2
  PIN pad_3_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 270 180 290 200 ;
    END
  END pad_3_2
  PIN connection_3_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 270 270 290 290 ;
    END
  END connection_3_3
  PIN pad_3_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 270 270 290 290 ;
    END
  END pad_3_3
  PIN connection_4_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 0 380 20 ;
    END
  END connection_4_0
  PIN pad_4_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 360 0 380 20 ;
    END
  END pad_4_0
  PIN connection_4_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 90 380 110 ;
    END
  END connection_4_1
  PIN pad_4_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 360 90 380 110 ;
    END
  END pad_4_1
  PIN connection_4_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 180 380 200 ;
    END
  END connection_4_2
  PIN pad_4_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 360 180 380 200 ;
    END
  END pad_4_2
  PIN connection_4_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 360 270 380 290 ;
    END
  END connection_4_3
  PIN pad_4_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 360 270 380 290 ;
    END
  END pad_4_3
  PIN connection_5_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 0 470 20 ;
    END
  END connection_5_0
  PIN pad_5_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 450 0 470 20 ;
    END
  END pad_5_0
  PIN connection_5_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 90 470 110 ;
    END
  END connection_5_1
  PIN pad_5_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 450 90 470 110 ;
    END
  END pad_5_1
  PIN connection_5_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 180 470 200 ;
    END
  END connection_5_2
  PIN pad_5_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 450 180 470 200 ;
    END
  END pad_5_2
  PIN connection_5_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 450 270 470 290 ;
    END
  END connection_5_3
  PIN pad_5_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 450 270 470 290 ;
    END
  END pad_5_3
  PIN connection_6_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 0 560 20 ;
    END
  END connection_6_0
  PIN pad_6_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 540 0 560 20 ;
    END
  END pad_6_0
  PIN connection_6_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 90 560 110 ;
    END
  END connection_6_1
  PIN pad_6_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 540 90 560 110 ;
    END
  END pad_6_1
  PIN connection_6_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 180 560 200 ;
    END
  END connection_6_2
  PIN pad_6_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 540 180 560 200 ;
    END
  END pad_6_2
  PIN connection_6_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 540 270 560 290 ;
    END
  END connection_6_3
  PIN pad_6_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 540 270 560 290 ;
    END
  END pad_6_3
  PIN connection_7_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 0 650 20 ;
    END
  END connection_7_0
  PIN pad_7_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 630 0 650 20 ;
    END
  END pad_7_0
  PIN connection_7_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 90 650 110 ;
    END
  END connection_7_1
  PIN pad_7_1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 630 90 650 110 ;
    END
  END pad_7_1
  PIN connection_7_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 180 650 200 ;
    END
  END connection_7_2
  PIN pad_7_2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 630 180 650 200 ;
    END
  END pad_7_2
  PIN connection_7_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 630 270 650 290 ;
    END
  END connection_7_3
  PIN pad_7_3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 630 270 650 290 ;
    END
  END pad_7_3
END interconnect_8x4

MACRO flush_hole_0
  CLASS PAD ;
  SIZE 40 BY 40 ;
  ORIGIN 0 0 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 0 20 40 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 20 0 40 40 ;
    END
  END pad
END flush_hole_0

MACRO pinhole_325px_met1
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met1 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 0 0 140 325 ;
    LAYER met2 ;
      RECT 0 0 140 325 ;
    LAYER met3 ;
      RECT 0 0 140 325 ;
    LAYER met4 ;
      RECT 0 0 140 325 ;
  END
END pinhole_325px_met1
MACRO pinhole_325px_met2
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met2 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 0 0 140 330 ;
    LAYER met2 ;
      RECT 0 0 140 330 ;
    LAYER met3 ;
      RECT 0 0 140 330 ;
    LAYER met4 ;
      RECT 0 0 140 330 ;
    LAYER met5 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met2

# Reminder to myself this is the previously working one
MACRO pinhole_325px_met3
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met3 ;
  SIZE 330 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 320 69 325 71 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 69 2 71 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 10 0 320 140 ;
    LAYER met2 ;
      RECT 10 0 320 140 ;
    LAYER met3 ;
      RECT 10 0 320 140 ;
    LAYER met4 ;
      RECT 10 0 320 140 ;
    LAYER met5 ;
      RECT 10 0 320 140 ;
    LAYER met6 ;
      RECT 10 0 320 140 ;
  END
END pinhole_325px_met3

# Reminder to myself this is the previously working one
MACRO pinhole_320px_0
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_0 ;
  SIZE 320 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300 60 320 80 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 0 60 20 80 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 20 0 300 140 ;
    LAYER met2 ;
      RECT 20 0 300 140 ;
    LAYER met3 ;
      RECT 20 0 300 140 ;
    LAYER met4 ;
      RECT 20 0 300 140 ;
    LAYER met5 ;
      RECT 20 0 300 140 ;
    LAYER met6 ;
      RECT 20 0 300 140 ;
  END
END pinhole_320px_0

MACRO pinhole_325px_met4
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met4 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 0 0 140 330 ;
    LAYER met2 ;
      RECT 0 0 140 330 ;
    LAYER met3 ;
      RECT 0 0 140 330 ;
    LAYER met4 ;
      RECT 0 0 140 330 ;
    LAYER met5 ;
      RECT 0 0 140 330 ;
    LAYER met6 ;
      RECT 0 0 140 330 ;
    LAYER met7 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met4
MACRO pinhole_325px_met5
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met5 ;
  SIZE 330 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310 60 330 80 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 0 60 20 80 ;
    END
  END pad
  OBS
    LAYER met1 ;
      RECT 20 0 310 140 ;
    LAYER met2 ;
      RECT 20 0 310 140 ;
    LAYER met3 ;
      RECT 20 0 310 140 ;
    LAYER met4 ;
      RECT 20 0 310 140 ;
    LAYER met5 ;
      RECT 20 0 310 140 ;
    LAYER met6 ;
      RECT 20 0 310 140 ;
    LAYER met7 ;
      RECT 20 0 310 140 ;
    LAYER met8 ;
      RECT 20 0 310 140 ;
    LAYER met9 ;
      RECT 20 0 310 140 ;
  END
END pinhole_325px_met5
MACRO pinhole_325px_met6
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met6 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met6 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met3 ;
      RECT 0 0 140 330 ;
    LAYER met4 ;
      RECT 0 0 140 330 ;
    LAYER met5 ;
      RECT 0 0 140 330 ;
    LAYER met6 ;
      RECT 0 0 140 330 ;
    LAYER met7 ;
      RECT 0 0 140 330 ;
    LAYER met8 ;
      RECT 0 0 140 330 ;
    LAYER met9 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met6
MACRO pinhole_325px_met7
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met7 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met7 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met4 ;
      RECT 0 0 140 330 ;
    LAYER met5 ;
      RECT 0 0 140 330 ;
    LAYER met6 ;
      RECT 0 0 140 330 ;
    LAYER met7 ;
      RECT 0 0 140 330 ;
    LAYER met8 ;
      RECT 0 0 140 330 ;
    LAYER met9 ;
      RECT 0 0 140 330 ;
    LAYER met10 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met7
MACRO pinhole_325px_met8
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met8 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met8 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met5 ;
      RECT 0 0 140 330 ;
    LAYER met6 ;
      RECT 0 0 140 330 ;
    LAYER met7 ;
      RECT 0 0 140 330 ;
    LAYER met8 ;
      RECT 0 0 140 330 ;
    LAYER met9 ;
      RECT 0 0 140 330 ;
    LAYER met10 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met8
MACRO pinhole_325px_met9
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met9 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met9 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met6 ;
      RECT 0 0 140 330 ;
    LAYER met7 ;
      RECT 0 0 140 330 ;
    LAYER met8 ;
      RECT 0 0 140 330 ;
    LAYER met9 ;
      RECT 0 0 140 330 ;
    LAYER met10 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met9

MACRO pinhole_325px_met10
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN pinhole_325px_met10 ;
  SIZE 140 BY 330 ;
  SYMMETRY X Y R90 ;
  PIN connection
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 325 71 327 ;
    END
  END connection
  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met10 ;
        RECT 69 0 71 2 ;
    END
  END pad
  OBS
    LAYER met7 ;
      RECT 0 0 140 330 ;
    LAYER met8 ;
      RECT 0 0 140 330 ;
    LAYER met9 ;
      RECT 0 0 140 330 ;
    LAYER met10 ;
      RECT 0 0 140 330 ;
  END
END pinhole_325px_met10

END LIBRARY
.,
