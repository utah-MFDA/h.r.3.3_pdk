

YPressurePump pr1         1  2   pressure=100k chemConcentration=100m
YPressurePump pr2         11 22  pressure=100k

Yserpentine_100px_0 serp1 1  3   2  4
Yserpentine_100px_0 serp2 11 13  22 24

Ydiffmix_25px_0 mix1      3  13  5  4  24 6

Yserpentine_100px_0 serp3 5  0  6  8
*Yserpentine_100px_0 serp3 5  100 6  8

*R1 8 0 1.0M

*Youtlet     out1  100 8

.tran 1m 10m 
.print tran V(1) V(3) V(4) V(6) V(8)
.end
