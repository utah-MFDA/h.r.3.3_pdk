

Vpp 1  0 PWL(0s 0V 3s 20V)
*Vpp 1  0 SIN(10V 20V 100Hz)

Vcc 11 0 0V

Yserpentine_100px_0  serp1 1  21 11 12

Ymembrane_cap_20px   mem1  22 31 capacitance=1n

Yserpentine_100px_0  serp2 32 0 12 13

* probe
Vpr1 31 32 0V 
Vpr2 21 22 0V

.tran 10ms 1s
.print tran V(22) V(31) I(Vpr1) I(Vpr2)
.end