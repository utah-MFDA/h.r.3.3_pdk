VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
END LIBRARY
