 
MACRO p_serpentine_0(L1.d, L2.d, turns.d)
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN p_serpentine_0 0 0 ;
  SIZE #L2*turns + 60# BY #L1 + 60# ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT #turns*L2+29.5# #((turns+1)%2)*L1+29.5# #turns*L2+30.5# #((turns+1)%2)*L1+30.5# ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 #L2*turns+60# #L1+60# ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END p_serpentine_0
