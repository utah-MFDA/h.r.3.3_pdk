

*Vpp 1  0 PWL(0s 0V 3s 20V)
Vpp 1  0 SIN(0V 10V 2meg)

Vcc 11 0 5V

Ychannel              serp1 1  21 11 12 length=100

Ymembrane_cap_20px    mem1  22 31 capacitance=1000u

Yserpentine_100px_0   serp2 32 0  12 13

* probe
Vpr1 31 32 0V 
Vpr2 22 21 0V

.tran 0.1ns 0.5us
.print tran V(22) V(31) V(1) I(Vpr1) I(Vpr2)
.end