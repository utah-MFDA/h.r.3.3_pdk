
*.options linsol type=klu

vs 1 0 PWL(0s 0kV 30ms 0kV 31ms 69kV 50ms 69kV 51ms 0V 1100.0ms 0V)

r1 22 21 1e11
Ymembrane_cap_20pxV_nlin_5_1 mem1 2 21 mem_r=540e-6 fl_ch_h=60e-6
*C_res=1e1


* probe sources
vp1 1 2 0V
vp2 0 22 0V

.tran 0.01ms 60ms 29ms 0.1ms
.print tran I(vp1) V(1) V(21)
.end
