

vs_f 1  0 0V

vs_p1 11 0 0
*PULSE(0kV 0   0.56   1m 1m 60m  300m)
vs_p2 12 0 PULSE(6.9kV 0   0.56   1m 1m 180m 300m)
vs_p3 13 0 0
*PULSE(0kV 0   0.68   1m 1m 120m 300m)

r1 1 2 1e11
r2 5 0 1e11


Yvalve_sw_20px_1_V              valv1 3 31 11 0  
Ymembrane_cap_20pxV_nlin_3_1 mem1  31 12 mem_r=504e-6 fl_ch_h=60e-6
Yvalve_sw_20px_1_V              valv2 31 4 13 0  

vp1 2 3 0V
vp2 4 5 0V 

.tran 0.008ms 2.1s 0.4s 0.01ms
.print tran I(vp1) I(vp2) V(11) V(12) V(13)
.end
