* serpentine 100 test

VC1 1 0 5V
VC2 2 0 8V
Yserpentine_100px_0 serp1 1 11 2 3
Yserpentine_100px_0 serp2 11 0 3 4 

.tran 1m 10m
.print tran I(vc1) V(3) V(11)
.end
