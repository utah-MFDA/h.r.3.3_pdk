

vs 1 0 PWL(0s 0V 5ms 0V 5.001ms 5V 10ms 5V)
r1 0 11 1k
r2 13 0 1k
Ymembrane_cap_20pxV_Pn mem1 2 1
*cap=1u

* probe sources
vp1 11 2 0V
vp2 2 13 0V

.tran 0.01ms 10ms
*.option post=2
.print tran I(vp2) I(vp1)
.end