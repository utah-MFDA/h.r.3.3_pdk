
MACRO serpentine_300px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN serpentine_300px_0 0 0 ;
  SIZE 420 BY 420 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 389.5 29.5 390.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 360 390 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END serpentine_300px_0
