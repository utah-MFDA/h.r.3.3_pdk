

YPressurePump prPump1 1 2   pressure=100k
YPressurePump prPump2 11 22 pressure=100k

Yserpentine_100px_0 serp1 1 3 2 4
Yserpentine_100px_0 serp2 11 13 22 24

Ydiffmix_25px_0 mix1 3 13 5 4 24 6

Yserpentine_100px_0 serp3 5 0 6 8

.tran 1m 10m 
.print tran V(1) V(3) V(5) V(8)
.end
