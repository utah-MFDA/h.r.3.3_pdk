*Test the channel objects

V1 1 0 5V 
Ychannel1 channel1 1 21
Ychannel1 channel2 22 0

V2 22 21 0V
* w=100u h=100u L=2m

.tran 1m 10m
.print tran I(v1)
.print tran I(v2)
.print tran V(1)
.print tran V(21)
.print tran V(22)
.end


