
MACRO pump_40px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_40px_0 0 0 ;
  SIZE 290 BY 135 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 69.5 30.5 70.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 259.5 69.5 260.5 70.5 ;
    END
  END out_fluid
  PIN a_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.5 29.5 75.5 30.5 ;
    END
  END a_in_air
  PIN a_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.5 109.5 75.5 110.5 ;
    END
  END a_out_air
  PIN b_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.5 29.5 145.5 30.5 ;
    END
  END b_in_air
  PIN b_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.5 109.5 145.5 110.5 ;
    END
  END b_out_air
  PIN c_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.5 29.5 215.5 30.5 ;
    END
  END c_in_air
  PIN c_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.5 109.5 215.5 110.5 ;
    END
  END c_out_air
  OBS
    LAYER met1 ;
      RECT 30 30 260 110 ;
    LAYER met2 ;
      RECT 30 30 260 110 ;
    LAYER met3 ;
      RECT 30 30 260 110 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_40px_0
