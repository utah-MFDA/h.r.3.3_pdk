*Test of the pump object

YPressurePump prpump 1 0

R1 1 0 50

.tran 1m 10m
.print tran V(1)
.end
