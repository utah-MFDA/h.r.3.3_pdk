*Test of the pump object

YEPressurePump prpump 1 0

R1 1 0 50

.tran 1m 10m
.print tran I(1)
.end
