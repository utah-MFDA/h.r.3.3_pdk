
MACRO optical_measure_100_5ch
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN optical_measure_100_5ch 0 0 ;
  SIZE 360 BY 120 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23 53 37 67 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 323 53 337 67 ;
    END
  END out_fluid
  OBS
    LAYER met1 ;
      RECT 30 30 330 90 ;
    LAYER met2 ;
      RECT 30 30 330 90 ;
    LAYER met3 ;
      RECT 40 30 320 90 ;
    LAYER met4 ;
      RECT 30 30 330 90 ;
    LAYER met5 ;
      RECT 40 30 320 90 ;
    LAYER met6 ;
      RECT 30 30 330 90 ;
    LAYER met7 ;
      RECT 30 30 330 90 ;
    LAYER met8 ;
      RECT 30 30 330 90 ;
    LAYER met9 ;
      RECT 30 30 330 90 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END optical_measure_100_5ch
