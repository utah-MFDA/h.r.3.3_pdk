* one stop valve per device

vs_f 1  0 0V

vs_p11 111 0 PULSE(69kV 0kV   0.56   5m 5m 60m  300m)
vs_p21 121 0 PULSE(69kV 0kV   0.56   5m 5m 180m 300m)
vs_p31 131 0 PULSE(69kV 0kV   0.68   5m 5m 120m 300m)

vs_p12 112 0 PULSE(69kV 0kV   0.56    5m 5m 60m  300m)
vs_p22 122 0 PULSE(69kV 0kV   0.56    5m 5m 180m 300m)
vs_p32 132 0 PULSE(69kV 0kV   0.68    5m 5m 120m 300m)

r1 1 2 1e11
r2 5 0 1e11


Yvalve_sw_20px_1_V              valv1 3  31 111 0 threshold_pressure_kPa=60e3 
Ymembrane_cap_20pxV_nlin_5_1 mem1  31 112 mem_r=540e-6 fl_ch_h=60e-6

Yvalve_sw_20px_1_V              valv2 31 32 121 0 threshold_pressure_kPa=60e3 
Ymembrane_cap_20pxV_nlin_5_1 mem2  32 122 mem_r=540e-6 fl_ch_h=60e-6

Yvalve_sw_20px_1_V              valv3 32 33 131 0 threshold_pressure_kPa=60e3 
Ymembrane_cap_20pxV_nlin_5_1 mem3  33 132 mem_r=540e-6 fl_ch_h=60e-6

vp1 2 3 0V
vp2 4 5 0V 

.tran 0.01ms 2.1s 0.4s 0.1ms
.print tran I(vp1) I(vp2) V(111) V(121) V(131)
.end
