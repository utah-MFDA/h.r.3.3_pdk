

vs 1 0 PWL(0s 0V 3ms 0V 3.001ms 5V 6ms 5V 6.001ms 0V 10ms 0V)
r1 1 2 1k
c1 3 0 1uF

vp 2 3 0V

.tran 0.01ms 10ms
*.option post=2
.print tran I(vs) I(vp)
.end