

MACRO p_serpentine_3(L1.d, L2.d, turns.d)
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN p_serpentine_3 0 0 ;
  SIZE #L2*turns + 60# BY #L1 + 60# ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END out_fluid
  OBS
    LAYER met2 ;
      RECT 30 30 #L2*turns+60# #L1+60# ;
    LAYER met3 ;
      RECT 30 30 #L2*turns+60# #L1+60# ;
    LAYER met4 ;
      RECT 30 30 #L2*turns+60# #L1+60# ;
    LAYER met5 ;
      RECT 30 30 #L2*turns+60# #L1+60# ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END p_serpentine_3
