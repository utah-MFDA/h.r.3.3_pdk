

YPressurePump prPump 1 2 pressure=100k

Yserpentine_100px_0 serp1 1 3 2 4
Yserpentine_100px_0 serp2 3 0 4 6
*Yserpentine_200px_0 serp3 5 0 6 0


.tran 1m 10m
.print tran V(1) V(6)
.end
