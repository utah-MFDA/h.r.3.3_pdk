
*.options linsol type=klu

vs 1 0 PWL(0s 0V 30ms 0V 40ms 500V 60ms 500V 70ms 0V 100.0ms 0V)

r1 0 21 1k
Ymembrane_cap_20pxV_nlin_4 mem1 2 21 mem_r=540e-6 fl_ch_h=60e-6
*C_res=1e1


* probe sources
vp1 1 2 0V

.tran 0.0001ms 100ms
.print tran I(vp1) V(1) V(2)
.end
