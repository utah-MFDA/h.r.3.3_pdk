*A simple rectangular channel

.hdl ./../../RectangularChannelElectrical.va
.options post=1
X1 1 0 RectangularChannelElectrical
VS 1 0 1
.dc VS 0 10 1
.end
