* serpentine 100 test


YPressurePump pr1  1  2   pressure=100k chemConcentration=100m

Ychannel serp1 1 11 2 3 length=10m
Ychannel serp2 11 0 3 4 length=10m
*c1 4 0 100u
*YOutput  out   4
*VCC 4 0 0V

*.preprocess addresistors nodcpath 1G
*.preprocess addresistors oneterminal 1G

.tran 1m 10m
.print tran V(3) V(11) 
*I(vcc)
.end
