

vs_f 1  0 5V
vs_p 11 0 PWL(0s 0V 3m 0v 3.1m 105kV 10m 015kV)

r1 1 2 1k
r2 5 0 1k
r3 11 12 1k
r4 13 0 1M

Yvalve_flow_20px_1 valv1 3 4 12 13   

vp1 2 3 0V
vp2 4 5 0V 

.tran 0.01 10ms
.print tran I(vp1) I(vp2)
.end